`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:29:39 07/12/2022 
// Design Name: 
// Module Name:    adder_IF 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder_IF(
    input [31:0] a1,
    output [31:0] b1
    );

assign b1= a1 +2'b01;




endmodule














